module adder_tb();

	logic [31:0] A, B, O;
	
	adder DUT(A, B, O);
	
	
	initial begin
	
	A = 32'b01000001001000000000000000000000; B = 32'b01000001001000000000000000000000; #10;
	assert (O === 32'b01000001101000000000000000000000) else $error("fail");
	
	A = 32'b01000001011100000000000000000000; B = 32'b11000001001000000000000000000000; #10;
	assert (O === 32'b01000000101000000000000000000000) else $error("fail");
	
	A = 32'b01000110010000001110010000000000; B = 32'b01000110101000000101100000000000; #10;
	assert (O === 32'b01000111000000000110010100000000) else $error("fail");
	
	
	end
	

endmodule

